module ExampleBlock();


endmodule
