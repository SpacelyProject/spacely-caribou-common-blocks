/fasic_home/lucahhot/Documents/spacely-caribou-common-blocks/spi_controller_interface/vivado/spi_controller_interface/spi_controller_interface.gen/sources_1/bd/spi_Sim/hdl/spi_Sim_wrapper.v