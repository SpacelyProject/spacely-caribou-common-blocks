module sp3_dual_rx();

   


   // Modules to add:
   // - lpgbtfpga-uplink
   // - sp3_demux
   // - cdc_rx
   // - mgt IP
   // - mgt IP reset synchronizer (?)




endmodule // sp3_dual_rx
