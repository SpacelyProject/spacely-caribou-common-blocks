//Remove Xilinx CDC IP for basic testing.
`define NO_CDC 1
module generic_spi_tb();


   //Controller signals
   logic [31:0] mem_write, mem_write_ptr, mem_read, mem_read_ptr;
   logic 	mem_write_strb, mem_write_ptr_reset, mem_read_strb, mem_read_ptr_reset;
   
   logic [31:0] transaction_count, transaction_len;
   logic 	master_spi_clk, poci, pico, cs_b, axi_clk, axi_resetn, run, spi_clk_gated, reset_b;
   logic [2:0] 	status;

   logic [31:0] loop_pattern, loop_iters, loop_counter;
   logic [7:0] 	loop_pattern_len;
   logic [2:0] 	loop_mode;
   
   
   generic_spi_controller controller (.*);

   
   //Peripheral spi_clk gets the spi_clk_gated output generated by the controller.
   logic 	spi_clk;
   
   assign spi_clk = spi_clk_gated;

   DUT_SP3 dut(.*);
   

   always begin
      #500;
      master_spi_clk = ~master_spi_clk;
   end

   always begin
      #10;
      axi_clk = ~axi_clk;

   end      
   				
   initial begin
      axi_clk = 0;
      master_spi_clk = 0;

      //Initial conditions: For Test 1, no loop.
      loop_mode = 0;
      loop_iters = 0;
      loop_pattern = 0;
      loop_pattern_len = 0;
      
      
      // Initial reset of both controller and peripheral.
      axi_resetn = 0;
      reset_b = 0;
      #10;
      axi_resetn = 1;
      reset_b = 1;
      

      // Wait at least one spi_clk period before starting.
      @(posedge master_spi_clk);
      @(posedge master_spi_clk);
      @(posedge master_spi_clk);
      

      // *********************************
      // * Test 1: Normal read/writeback *
      // *********************************

      // Write 10101010 to the address 00_1000_0000
      // Remember that the memory is little-endian! bit [0] is
      // transmitted first.
  
      @(posedge axi_clk) ;
      mem_write_strb = 1'b1;
      mem_write = 32'b01010101_0000_0001_00_1;
      @(posedge axi_clk) ;
      mem_write_strb = 1'b0;
      transaction_len = 19;
      @(posedge axi_clk);
      
      do_transaction();
      

      // Now read the stame address. Remember to reset the mem_write_ptr
      @(posedge axi_clk) ;
      mem_write_ptr_reset = 1'b1;
      @(posedge axi_clk) ;
      mem_write_ptr_reset = 1'b0;
      mem_write_strb = 1'b1;
      mem_write = 32'b00000000_0000_0001_00_0;
      @(posedge axi_clk) ;
      mem_write_strb = 1'b0;
      transaction_len = 20;

      do_transaction();

      //Remember that the first 12 bits of any read will be garbage.
      //1b offset + 1b WnR + 10b address.
      $display("mem_read: %b",mem_read[19:12]);
      if(mem_read[19:12] == 8'b01010101)
	$display("Test 1 -- SUCCESS!");
      else
	$display("Test 1 -- FAIL");
      
      
      // **********************************
      // * Test 2: Normal Config Chain Push *
      // **********************************
      //Push a miscellaneous clock-like pattern into the config chain.
       @(posedge axi_clk) ;
      mem_write_ptr_reset = 1'b1;
      @(posedge axi_clk) ;
      mem_write_ptr_reset = 1'b0;

      //Recall that to mimic a real AXI interface, mem_write_strb
      //gets asserted one clock cycle earlier than the data actually arrives.
      mem_write_strb = 1'b1;
      @(posedge axi_clk);
      mem_write = 32'b011011011011011011011_1000_0000_01_1;
      @(posedge axi_clk) ;
      mem_write_strb = 1'b0;
      mem_write = 32'b11001100110011001100110011001100;
       @(posedge axi_clk) ;
     // mem_write_strb = 1'b0;
      transaction_len = 64;

      do_transaction();
      

      // **********************************
      // * Test 3: Loop Config Chain Push *
      // **********************************
      //20 x 10b = twice through the 100-bit config chain.
       @(posedge axi_clk) ;
      mem_write_ptr_reset = 1'b1;
      @(posedge axi_clk) ;
      mem_write_ptr_reset = 1'b0;
      mem_write_strb = 1'b1;
      mem_write = 32'b1000_0000_01_1;
       @(posedge axi_clk) ;
      mem_write_strb = 1'b0;
      transaction_len = 11;
      @(posedge axi_clk) ;
      loop_mode = 1;
      @(posedge axi_clk) ;
      loop_pattern = 32'b0111011010;
      @(posedge axi_clk) ;
      loop_pattern_len = 10;
      @(posedge axi_clk) ;
      loop_iters = 20;
      @(posedge axi_clk);


      do_transaction();
      
		     

      
      $finish();
      


   end // initial begin

   task do_transaction();
      //Send transaction
      @(posedge axi_clk);
      run = 1;
      @(posedge axi_clk);
      run = 0;
      
      // Wait for transaction to complete
      while(status > 0) @(posedge axi_clk);

      // Wait for one more posedge of spi_clk to allow the ASIC state
      // machine to reset.  
      @(posedge spi_clk_gated);
      


   endtask // do_transaction

     initial begin
      $dumpfile("DB.vcd");
      $dumpvars(0, generic_spi_tb); //Dump variables from level 0 and up 
   end
   

endmodule // generic_spi_tb


